`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:25:05 12/28/2020 
// Design Name: 
// Module Name:    pacman_behavior 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module pacman_behavior(input wire [9:0] pacx,
								input wire [8:0] pacy,
								input wire [9:0] ghostx,
								input wire [8:0] ghosty,
								
    );


endmodule
